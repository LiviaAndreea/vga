module ClkDivider (

    input EN,
	 input clock_div,
    output clk,
    input rst
 );
    


 endmodule

 






